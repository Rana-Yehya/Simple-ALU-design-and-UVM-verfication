package ALU_pkg;
  import uvm_pkg::*;
	`include "uvm_macros.svh"
  	`include "ALU_sequencer.sv"
	`include "ALU_monitor.sv"
	`include "ALU_driver.sv"
	`include "ALU_agent.sv"
	`include "ALU_scoreboard.sv"
	`include "ALU_config.sv"
	`include "ALU_env.sv"
	`include "ALU_test.sv"
	`include "ALU_coverage.sv"
endpackage: ALU_pkg
